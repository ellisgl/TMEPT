`timescale 1ns / 1ps
`default_nettype none
////////////////////////////////////////////////////////////////////////////////
// ROM Module
// 32k x 8-bit Read-Only Memory initialized from external hex file.
////////////////////////////////////////////////////////////////////////////////
module rom (
    input  wire [14:0] ADDR, // 15-bit
    input  wire        CS,   // active high
    output wire  [7:0] DO    // 8-bit
);

    reg [7:0] rom [0:32767]; // 32kbyte ROM space.

    // Initialize ROM from the Intel hex memory file generated by the build.

    initial $readmemh("build/tmept.mem", rom, 0, 32767);

    // Output ROM value if chip selected. If not chip selected, output high impedance.
    assign DO = CS ? rom[ADDR] : 8'bzzzzzzzz;
endmodule
`default_nettype wire
